library IEEE;
use IEEE.std_logic_1164.all;

package register_array_typev2 is
  type registerArray is array(0 to 7) of std_logic;
end package register_array_typev2;